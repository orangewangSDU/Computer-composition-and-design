library verilog;
use verilog.vl_types.all;
entity multiply_vlg_check_tst is
    port(
        qq0             : in     vl_logic;
        qq1             : in     vl_logic;
        qq2             : in     vl_logic;
        qq3             : in     vl_logic;
        qq4             : in     vl_logic;
        qq5             : in     vl_logic;
        qq6             : in     vl_logic;
        qq7             : in     vl_logic;
        qq8             : in     vl_logic;
        qq9             : in     vl_logic;
        qq10            : in     vl_logic;
        qq11            : in     vl_logic;
        qq12            : in     vl_logic;
        qq13            : in     vl_logic;
        qq14            : in     vl_logic;
        qq15            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end multiply_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity multiply_vlg_vec_tst is
end multiply_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity multiply is
    port(
        qq7             : out    vl_logic;
        A0              : in     vl_logic;
        B0              : in     vl_logic;
        B1              : in     vl_logic;
        A1              : in     vl_logic;
        B2              : in     vl_logic;
        A2              : in     vl_logic;
        B3              : in     vl_logic;
        A3              : in     vl_logic;
        B4              : in     vl_logic;
        A4              : in     vl_logic;
        B5              : in     vl_logic;
        A5              : in     vl_logic;
        B6              : in     vl_logic;
        A6              : in     vl_logic;
        B7              : in     vl_logic;
        A7              : in     vl_logic;
        qq6             : out    vl_logic;
        qq5             : out    vl_logic;
        qq4             : out    vl_logic;
        qq3             : out    vl_logic;
        qq2             : out    vl_logic;
        qq1             : out    vl_logic;
        qq0             : out    vl_logic;
        qq15            : out    vl_logic;
        qq14            : out    vl_logic;
        qq13            : out    vl_logic;
        qq12            : out    vl_logic;
        qq11            : out    vl_logic;
        qq10            : out    vl_logic;
        qq9             : out    vl_logic;
        qq8             : out    vl_logic
    );
end multiply;

library verilog;
use verilog.vl_types.all;
entity ex1_vlg_vec_tst is
end ex1_vlg_vec_tst;
